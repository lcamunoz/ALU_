library verilog;
use verilog.vl_types.all;
entity ALU_final_vlg_vec_tst is
end ALU_final_vlg_vec_tst;
